package comm_pkg;

endpackage